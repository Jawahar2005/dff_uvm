interface dff_interface;
  //Paramater 
  parameter WIDTH = 4;
 
  logic clk,rst;
  logic [WIDTH-1:0] din;
  logic [WIDTH-1:0] dout;
  
endinterface
